-- Computer Architecture - Technical University of Crete
-- Speculative Tomasulo’s Algorithm
-- N. Kyparissas, A. Kampylafkas

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ROB IS
PORT (
	CLK : IN STD_LOGIC;
	RST : IN STD_LOGIC;
	-- ISSUE
	PC : IN STD_LOGIC_VECTOR(9 DOWNTO 0); -- HERE: OUR PC COUNTER
	ISSUE_WE : IN STD_LOGIC;
	INSTRUCTION : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
	Q_FOR_NEW_INSTR : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); -- = TAIL 
	-- NEW INSTRUCTION
	Q_RS_ROB : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); -- IN CASE THE DATA YOU'VE BEEN ASKING IN REGISTER FILE IS NOT VALID
	Q_RT_ROB : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	DATA_RS_ROB : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	DATA_RT_ROB : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	DATA_RS_ROB_VALID : OUT STD_LOGIC;
	DATA_RT_ROB_VALID : OUT STD_LOGIC;
	-- CDB
	CDB_V : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	CDB_Q : IN STD_LOGIC_VECTOR(3 DOWNTO 0); 
	-- RF (COMMIT)
	ROB_VALUE : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	ROB_RD : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
	RF_WE : OUT STD_LOGIC;
	-- EXCEPTION
	EXCEPTION_PC : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
	EXCEPTION_ROB_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); 
	EXCEPTION_FLAG : IN STD_LOGIC; 
	EXCEPTION_ROB_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0)); -- INTERNAL EXCEPTION - SOME FU SENDS BACK THIS ROB, IF NOT, WE CAN EASILY GET THAT FROM PC NUMBER
END ROB;

ARCHITECTURE BEHAVIORAL OF ROB IS
	SIGNAL TAIL, HEAD : UNSIGNED(3 DOWNTO 0) := (OTHERS => '0');
	SIGNAL EXCEPTION_ROB_OUT_SIG : STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '1');
	
	-- 4B (51 DOWNTO 48): INSTRUCTION, 10B (47 DOWNTO 38): PC, 5B (37 DOWNTO 33): RD, 32B (32 DOWNTO 1): VALUE, 1B (0): DONE
	TYPE ROB_REGISTER IS ARRAY(14 DOWNTO 0) OF STD_LOGIC_VECTOR(51 DOWNTO 0);
	SIGNAL ROB_REG : ROB_REGISTER := (OTHERS => (OTHERS => '0'));

BEGIN

	PROCESS
	BEGIN

		WAIT UNTIL RISING_EDGE(CLK);

		IF (RST = '1') THEN
			-- RF
			RF_WE <= '0';
			ROB_VALUE <= (OTHERS => '0');
			ROB_RD <= (OTHERS => '0');
			-- NEW INSTRUCTION
			Q_RS_ROB <= (OTHERS => '1');
			Q_RT_ROB <= (OTHERS => '1');
			DATA_RS_ROB <= (OTHERS => '0');
			DATA_RT_ROB <= (OTHERS => '0');
			DATA_RS_ROB_VALID <= '0';
			DATA_RT_ROB_VALID <= '0';
			-- EXCEPTION
			EXCEPTION_PC <= (OTHERS => '0');
			EXCEPTION_ROB_OUT_SIG <= (OTHERS => '1'); -- "1111" MEANS THERE IS NO EXCEPTION
			-- INTERNAL ROB SIGNALS
			TAIL <= (OTHERS => '0');
			HEAD <= (OTHERS => '0');
			ROB_REG <= (OTHERS => (OTHERS => '0'));
		ELSE
			IF EXCEPTION_FLAG = '1' THEN

				EXCEPTION_PC <= ROB_REG(TO_INTEGER(UNSIGNED(EXCEPTION_ROB_IN)))(47 DOWNTO 38); -- PC
				EXCEPTION_ROB_OUT_SIG <= EXCEPTION_ROB_IN; 

				-- FLUSHING ROB REGISTRIES
				IF UNSIGNED(EXCEPTION_ROB_IN) <= TAIL THEN 
					-- L_0: FOR I IN TO_INTEGER(UNSIGNED(EXCEPTION_ROB_IN)) TO TO_INTEGER(TAIL-1) LOOP -- THIS LINE IS NOT SYNTHESIZABLE, REPLACED BY THE TWO LINES BELOW
					L_0: FOR I IN 0 TO 14 LOOP
						IF I >= TO_INTEGER(UNSIGNED(EXCEPTION_ROB_IN)) AND I <= TO_INTEGER(TAIL-1) THEN
							ROB_REG(I) <= (OTHERS => '0');            
						END IF;
					END LOOP L_0;   
				ELSE 
					-- L_1: FOR I IN TO_INTEGER(UNSIGNED(EXCEPTION_ROB_IN)) TO 14 LOOP -- THIS LINE IS NOT SYNTHESIZABLE, REPLACED BY THE TWO LINES BELOW
					L_1: FOR I IN 0 TO 14 LOOP
						IF I >= TO_INTEGER(UNSIGNED(EXCEPTION_ROB_IN)) THEN
							ROB_REG(I) <= (OTHERS => '0');            
						END IF;
					END LOOP L_1;
					-- L_2: FOR I IN 0 TO TO_INTEGER(TAIL-1) LOOP -- THIS LINE IS NOT SYNTHESIZABLE, REPLACED BY THE TWO LINES BELOW
					L_2: FOR I IN 0 TO 14 LOOP
						IF I <= TO_INTEGER(TAIL-1) THEN 
							ROB_REG(I) <= (OTHERS => '0'); 
						END IF;           
					END LOOP L_2;
				END IF;           
			ELSE
				-- WE DON'T HAVE AN EXCEPTION (ANY MORE? ;) ), RESET EXCEPTION ROB
				IF EXCEPTION_ROB_OUT_SIG /= "1111" THEN
					TAIL <= UNSIGNED(EXCEPTION_ROB_IN); -- TAIL VALUE NEEDS TO BE UPDATED AFTER THE EXCEPTION, SO THAT THE RESERVATION STATIONS WONT DELETE THE WRONG VALUES
					EXCEPTION_ROB_OUT_SIG <= (OTHERS => '1'); 
				END IF;

				IF CDB_Q /= "1111" THEN -- CDB IS BROADCASTING SOMETHING
					ROB_REG(TO_INTEGER(UNSIGNED(CDB_Q)))(32 DOWNTO 1) <= CDB_V;
					ROB_REG(TO_INTEGER(UNSIGNED(CDB_Q)))(0) <= '1';
				END IF;

				-- COMMIT
				IF ROB_REG(TO_INTEGER(HEAD))(0) = '1' THEN 
					ROB_VALUE <= ROB_REG(TO_INTEGER(HEAD))(32 DOWNTO 1);
					ROB_RD <= ROB_REG(TO_INTEGER(HEAD))(37 DOWNTO 33);
					RF_WE <= '1';
					ROB_REG(TO_INTEGER(HEAD)) <= (OTHERS => '0'); -- FLUSHING ROB REGISTRY
					IF HEAD = 14 THEN
						HEAD <= (OTHERS => '0'); -- "1111" NOT ALLOWED!
					ELSE 
						HEAD <= HEAD + 1;
					END IF;
				ELSIF TO_INTEGER(UNSIGNED(CDB_Q)) = HEAD THEN -- CDB_Q = HEAD: WRITE-FIRST, ESSENTIAL FOR CORNER CASES (SIMULTANEOUS ISSUE RS/RT, CDB BROADCAST)
					ROB_VALUE <= CDB_V;
					ROB_RD <= ROB_REG(TO_INTEGER(HEAD))(37 DOWNTO 33);
					RF_WE <= '1';
					ROB_REG(TO_INTEGER(HEAD)) <= (OTHERS => '0'); -- FLUSHING ROB REGISTRY
					IF HEAD = 14 THEN
						HEAD <= (OTHERS => '0'); -- "1111" NOT ALLOWED!
					ELSE 
						HEAD <= HEAD + 1;
					END IF;
				ELSE    
					RF_WE <= '0';
				END IF;

				-- NEW INSTRUCTION ISSUE
				-- TAIL ALWAYS SHOWS THE ROB TO BE OCCUPIED BY THE NEXT INSTRUCTION
				IF ISSUE_WE = '1' THEN
					ROB_REG(TO_INTEGER(TAIL))(51 DOWNTO 48) <= INSTRUCTION(18 DOWNTO 15); -- WHAT KIND OF INSTR?
					ROB_REG(TO_INTEGER(TAIL))(47 DOWNTO 38) <= PC; -- PC
					ROB_REG(TO_INTEGER(TAIL))(37 DOWNTO 33) <= INSTRUCTION(14 DOWNTO 10); -- RD
					ROB_REG(TO_INTEGER(TAIL))(0) <= '0'; -- DONE
					IF TAIL = 14 THEN
						TAIL <= (OTHERS => '0'); -- "1111" NOT ALLOWED!
					ELSE 
						TAIL <= TAIL + 1;
					END IF;
				END IF;

				-- NEW INSTRUCTION ASKS FOR RS AND RT:
				Q_RS_ROB <= "1111"; -- INSTRUCTION'S RS OR RT NOT FOUND YET	
				Q_RT_ROB <= "1111";
				DATA_RS_ROB_VALID <= '0';
				DATA_RT_ROB_VALID <= '0';
				-- IF THE SEARCHES BELOW DONT FIND ANYTHING, Q_RS_ROB AND Q_RT_ROB VALUES WILL REMAIN "1111"
				-- SO THAT RESERVATION STATIONS WILL NEGLECT ROB AND LOAD DATA FROM RF
				IF CDB_Q /= "1111" AND ROB_REG(TO_INTEGER(UNSIGNED(CDB_Q)))(37 DOWNTO 33) = INSTRUCTION(9 DOWNTO 5) THEN -- IF CDB IS BROACASTING A VALUE FOR INSTRUCTION'S RS
					Q_RS_ROB <= CDB_Q; -- Q
					DATA_RS_ROB <= CDB_V; -- VALUE
					DATA_RS_ROB_VALID <= '1'; -- VALID
				ELSIF CDB_Q /= "1111" AND ROB_REG(TO_INTEGER(UNSIGNED(CDB_Q)))(37 DOWNTO 33) = INSTRUCTION(4 DOWNTO 0) THEN -- IF CDB IS BROACASTING A VALUE FOR INSTRUCTION'S RT
					Q_RT_ROB <= CDB_Q; -- Q
					DATA_RT_ROB <= CDB_V; -- VALUE
					DATA_RT_ROB_VALID <= '1'; -- VALID
				ELSIF HEAD < TAIL THEN -- IF CDB IS NOT BROACASTING ANYTHING RELEVANT, LOOK FOR THE MOST RECENT VALUE STORED IN ROB FOR INSTRUCTION'S RS AND RT
					-- L_3: FOR I IN TO_INTEGER(HEAD) TO TO_INTEGER(TAIL-1) LOOP -- THIS LINE IS NOT SYNTHESIZABLE, REPLACED BY THE TWO LINES BELOW
					L_3: FOR I IN 0 TO 14 LOOP
						IF I >= TO_INTEGER(HEAD) AND I <= TO_INTEGER(TAIL-1) THEN	
							-- RS
							IF ROB_REG(I)(37 DOWNTO 33) = INSTRUCTION(9 DOWNTO 5) THEN -- IF ROB'S RD = INSTRUCTION'S RS
								Q_RS_ROB <= STD_LOGIC_VECTOR(TO_UNSIGNED(I, Q_RS_ROB'LENGTH)); -- Q
								DATA_RS_ROB <= ROB_REG(I)(32 DOWNTO 1); -- VALUE
								DATA_RS_ROB_VALID <= ROB_REG(I)(0); -- VALID OR NOT
							END IF;
							-- RT
							IF ROB_REG(I)(37 DOWNTO 33) = INSTRUCTION(4 DOWNTO 0) THEN -- IF ROB'S RD = INSTRUCTION'S RT
								Q_RT_ROB <= STD_LOGIC_VECTOR(TO_UNSIGNED(I, Q_RT_ROB'LENGTH)); -- Q
								DATA_RT_ROB <= ROB_REG(I)(32 DOWNTO 1); -- VALUE
								DATA_RT_ROB_VALID <= ROB_REG(I)(0); -- VALID OR NOT
							END IF;
						END IF;
					END LOOP L_3;    
				ELSIF HEAD /= TAIL THEN 
					-- HEAD TO END
					-- L_4: FOR I IN TO_INTEGER(HEAD) TO 14 LOOP -- THIS LINE IS NOT SYNTHESIZABLE, REPLACED BY THE TWO LINES BELOW
					L_4: FOR I IN 0 TO 14 LOOP   
						IF I >= TO_INTEGER(HEAD) THEN
							-- RS
							IF ROB_REG(I)(37 DOWNTO 33) = INSTRUCTION(9 DOWNTO 5) THEN -- IF ROB'S RD = INSTRUCTION'S RS
								Q_RS_ROB <= STD_LOGIC_VECTOR(TO_UNSIGNED(I, Q_RS_ROB'LENGTH)); -- Q
								DATA_RS_ROB <= ROB_REG(I)(32 DOWNTO 1); -- VALUE
								DATA_RS_ROB_VALID <= ROB_REG(I)(0); -- VALID OR NOT
							END IF;
							-- RT
							IF ROB_REG(I)(37 DOWNTO 33) = INSTRUCTION(4 DOWNTO 0) THEN -- IF ROB'S RD = INSTRUCTION'S RT
								Q_RT_ROB <= STD_LOGIC_VECTOR(TO_UNSIGNED(I, Q_RT_ROB'LENGTH));-- Q
								DATA_RT_ROB <= ROB_REG(I)(32 DOWNTO 1); -- VALUE
								DATA_RT_ROB_VALID <= ROB_REG(I)(0); -- VALID OR NOT
							END IF;     
						END IF;      
					END LOOP L_4;
					-- END TO TAIL
					-- L_5: FOR I IN 0 TO TO_INTEGER(TAIL-1) LOOP -- THIS LINE IS NOT SYNTHESIZABLE, REPLACED BY THE TWO LINES BELOW
					L_5: FOR I IN 0 TO 14 LOOP
						IF I <= TO_INTEGER(TAIL-1) THEN
							-- RS
							IF ROB_REG(I)(37 DOWNTO 33) = INSTRUCTION(9 DOWNTO 5) THEN -- IF ROB'S RD = INSTRUCTION'S RS
								Q_RS_ROB <= STD_LOGIC_VECTOR(TO_UNSIGNED(I, Q_RS_ROB'LENGTH)); -- Q
								DATA_RS_ROB <= ROB_REG(I)(32 DOWNTO 1); -- VALUE
								DATA_RS_ROB_VALID <= ROB_REG(I)(0); -- VALID OR NOT
							END IF;
							-- RT
							IF ROB_REG(I)(37 DOWNTO 33) = INSTRUCTION(4 DOWNTO 0) THEN -- IF ROB'S RD = INSTRUCTION'S RT
								Q_RT_ROB <= STD_LOGIC_VECTOR(TO_UNSIGNED(I, Q_RT_ROB'LENGTH)); -- Q
								DATA_RT_ROB <= ROB_REG(I)(32 DOWNTO 1); -- VALUE
								DATA_RT_ROB_VALID <= ROB_REG(I)(0); -- VALID OR NOT
							END IF;     
						END IF;       
					END LOOP L_5;
				END IF;   
			END IF;
		END IF;
	END PROCESS;

	-- TAIL ALWAYS SHOWS THE ROB TO BE OCCUPIED BY THE NEXT INSTRUCTION
	Q_FOR_NEW_INSTR <= STD_LOGIC_VECTOR(TAIL);
	EXCEPTION_ROB_OUT <= EXCEPTION_ROB_OUT_SIG;

END BEHAVIORAL;
