-- COMPUTER ARCHITECTURE - TECHNICAL UNIVERSITY OF CRETE
-- SPECULATIVE TOMASULO’S ALGORITHM
-- N. KYPARISSAS, A. KAMPYLAFKAS

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY RESERVATION_STATIONS_ARITH IS
	PORT(
		CLK : IN STD_LOGIC;
		RST : IN STD_LOGIC;
		-- ISSUE SIGNALS
		INSTRUCTION : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
		ACK : OUT STD_LOGIC; -- LETTING ISSUE STG KNOW THAT THIS RS IS ACCEPTING ITS CURRENT INSTR
		-- ROB SIGNALS
		Q_RS_ROB : IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- IN CASE THE DATA YOU'VE BEEN ASKING IN REGISTER FILE IS NOT VALID
		Q_RT_ROB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		DATA_RS_ROB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_RT_ROB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_RS_ROB_VALID : IN STD_LOGIC;
		DATA_RT_ROB_VALID : IN STD_LOGIC;
		Q_FOR_NEW_INSTR : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		EXCEPTION_ROB : IN STD_LOGIC_VECTOR(3 DOWNTO 0); 
		-- RF SIGNALS
		DATA_RS_RF : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_RT_RF : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		-- FU SIGNALS
		FU_Q : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);  
		FU_V1 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		FU_V2 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		FU_OP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		-- CDB SIGNALS
		CDB_Q : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CDB_V : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		CDB_Q_ACCESS_GRANTED : IN STD_LOGIC_VECTOR (1 DOWNTO 0)); -- EVERY TIME WE SEND A VALUE TO BE COMPUTED, WE COUNT UP UNTIL THE PIPELINE IS FULL.
		-- EVERY TIME CDB TAKES A VALUE, WE COUNT DOWN AND THAT MEANS WE CAN SEND ANOTHER VALUE. 
END RESERVATION_STATIONS_ARITH;

ARCHITECTURE BEHAVIORAL OF RESERVATION_STATIONS_ARITH IS
	-- (78 DOWNTO 75): ROB TAG, (74): BUSY, (73 DOWNTO 72): OP, (71 DOWNTO 40): V1 , (39 DOWNTO 36): Q1, (35 DOWNTO 4): V2, (3 DOWNTO 0): Q2
	TYPE RESERVATION_STATIONS IS ARRAY(2 DOWNTO 0) OF STD_LOGIC_VECTOR(78 DOWNTO 0); -- ARITHMETIC FU HAS 3 RESERVATION STATIONS
	SIGNAL RESERVATION_STATION : RESERVATION_STATIONS := (OTHERS => (OTHERS => '0'));	
	SIGNAL COUNTER : UNSIGNED(1 DOWNTO 0) := (OTHERS => '0');
	SIGNAL RS0_WAIT_FOR_RF, RS1_WAIT_FOR_RF, RS2_WAIT_FOR_RF, ACK_SIG : STD_LOGIC := '0';
	
BEGIN

	PROCESS
	BEGIN
	
		WAIT UNTIL RISING_EDGE(CLK);
		
		IF (RST = '1') THEN
			RESERVATION_STATION <= (OTHERS => (OTHERS => '0'));
			FU_Q <= "1111"; -- THERE IS NO SUCH RS, WE ARE SENDING OUT NOTHING
			FU_V1 <= (OTHERS => '0');
			FU_V2 <= (OTHERS => '0');
			FU_OP <= (OTHERS => '0');
			COUNTER <= (OTHERS => '0');
			RS0_WAIT_FOR_RF <= '0';
			RS1_WAIT_FOR_RF <= '0';
			RS2_WAIT_FOR_RF <= '0';
		-- EXCEPTION DETECTED BY ROB: KAZANAKI (FLUSHING)
		ELSIF EXCEPTION_ROB /= "1111" THEN	
			-- FLUSHING ROB REGISTRIES
			IF UNSIGNED(EXCEPTION_ROB) < UNSIGNED(Q_FOR_NEW_INSTR) THEN 
				-- L_1: FOR I IN TO_INTEGER(UNSIGNED(EXCEPTION_ROB)) TO TO_INTEGER(UNSIGNED(Q_FOR_NEW_INSTR))-1 LOOP -- THIS LINE IS NOT SYNTHESIZABLE, REPLACED BY THE TWO LINES BELOW
				L_1: FOR I IN 0 TO 14 LOOP 
					IF I >= TO_INTEGER(UNSIGNED(EXCEPTION_ROB)) AND I <= TO_INTEGER(UNSIGNED(Q_FOR_NEW_INSTR))-1 THEN    
						IF TO_INTEGER(UNSIGNED(RESERVATION_STATION(0)(78 DOWNTO 75))) = I THEN -- IF THE RS' TAG IS NEWER THAN THE EXCEPTION
							RESERVATION_STATION(0) <= (OTHERS => '0'); -- FLUSH IT
						END IF;
						IF TO_INTEGER(UNSIGNED(RESERVATION_STATION(1)(78 DOWNTO 75))) = I THEN -- IF THE RS' TAG IS NEWER THAN THE EXCEPTION
							RESERVATION_STATION(1) <= (OTHERS => '0'); -- FLUSH IT
						END IF;
						IF TO_INTEGER(UNSIGNED(RESERVATION_STATION(2)(78 DOWNTO 75))) = I THEN -- IF THE RS' TAG IS NEWER THAN THE EXCEPTION
							RESERVATION_STATION(2) <= (OTHERS => '0'); -- FLUSH IT
						END IF;
					END IF;
				END LOOP L_1;    
			ELSE 
				-- L_2: FOR I IN TO_INTEGER(UNSIGNED(EXCEPTION_ROB)) TO 14 LOOP -- THIS LINE IS NOT SYNTHESIZABLE, REPLACED BY THE TWO LINES BELOW
				L_2: FOR I IN 0 TO 14 LOOP
					IF I >= TO_INTEGER(UNSIGNED(EXCEPTION_ROB)) THEN
						IF TO_INTEGER(UNSIGNED(RESERVATION_STATION(0)(78 DOWNTO 75))) = I THEN -- IF THE RS' TAG IS NEWER THAN THE EXCEPTION
							RESERVATION_STATION(0) <= (OTHERS => '0'); -- FLUSH IT
						END IF;
						IF TO_INTEGER(UNSIGNED(RESERVATION_STATION(1)(78 DOWNTO 75))) = I THEN -- IF THE RS' TAG IS NEWER THAN THE EXCEPTION
							RESERVATION_STATION(1) <= (OTHERS => '0'); -- FLUSH IT
						END IF;
						IF TO_INTEGER(UNSIGNED(RESERVATION_STATION(2)(78 DOWNTO 75))) = I THEN -- IF THE RS' TAG IS NEWER THAN THE EXCEPTION
							RESERVATION_STATION(2) <= (OTHERS => '0'); -- FLUSH IT
						END IF;
					END IF;
				END LOOP L_2;
				-- L_3: FOR I IN 0 TO TO_INTEGER(UNSIGNED(Q_FOR_NEW_INSTR))-1 LOOP -- THIS LINE IS NOT SYNTHESIZABLE, REPLACED BY THE TWO LINES BELOW
				L_3: FOR I IN 0 TO 14 LOOP
					IF I <= TO_INTEGER(UNSIGNED(Q_FOR_NEW_INSTR))-1 THEN
						IF TO_INTEGER(UNSIGNED(RESERVATION_STATION(0)(78 DOWNTO 75))) = I THEN -- IF THE RS' TAG IS NEWER THAN THE EXCEPTION
							RESERVATION_STATION(0) <= (OTHERS => '0'); -- FLUSH IT
						END IF;
						IF TO_INTEGER(UNSIGNED(RESERVATION_STATION(1)(78 DOWNTO 75))) = I THEN -- IF THE RS' TAG IS NEWER THAN THE EXCEPTION
							RESERVATION_STATION(1) <= (OTHERS => '0'); -- FLUSH IT
						END IF;
						IF TO_INTEGER(UNSIGNED(RESERVATION_STATION(2)(78 DOWNTO 75))) = I THEN -- IF THE RS' TAG IS NEWER THAN THE EXCEPTION
							RESERVATION_STATION(2) <= (OTHERS => '0'); -- FLUSH IT
						END IF;
					END IF;
				END LOOP L_3;
			END IF;       
		ELSE
			-- ACCEPTING (OR NOT) AN ISSUED INSTRUCTION
			IF INSTRUCTION(18 DOWNTO 17) = "01" AND ACK_SIG = '1' THEN -- IF THE INSTRUCTION IS AN ARITHMETIC ONE AND THERE IS AN AVAILABLE RS
				IF RESERVATION_STATION(0)(74) = '0' THEN -- IF RS(0) AVAILABLE WRITE HERE ELSE KEEP SEARCHING FOR AVAILABLE RS
					RESERVATION_STATION(0)(74) <= '1';
					RESERVATION_STATION(0)(73 DOWNTO 72) <= INSTRUCTION(16 DOWNTO 15); -- FOP
					RESERVATION_STATION(0)(78 DOWNTO 75) <= Q_FOR_NEW_INSTR; -- TAG FROM ROB
					RS0_WAIT_FOR_RF <= '1'; -- FILL RS FROM RF IN THE NEXT CYCLE
				ELSIF RESERVATION_STATION(1)(74) = '0' THEN
					RESERVATION_STATION(1)(74) <= '1';
					RESERVATION_STATION(1)(73 DOWNTO 72) <= INSTRUCTION(16 DOWNTO 15); -- FOP
					RESERVATION_STATION(1)(78 DOWNTO 75) <= Q_FOR_NEW_INSTR; -- TAG FROM ROB
					RS1_WAIT_FOR_RF <= '1'; -- FILL RS FROM RF IN THE NEXT CYCLE
				ELSIF RESERVATION_STATION(2)(74) = '0' THEN
					RESERVATION_STATION(2)(74) <= '1';
					RESERVATION_STATION(2)(73 DOWNTO 72) <= INSTRUCTION(16 DOWNTO 15); -- FOP
					RESERVATION_STATION(2)(78 DOWNTO 75) <= Q_FOR_NEW_INSTR; -- TAG FROM ROB
					RS2_WAIT_FOR_RF <= '1'; -- FILL RS FROM RF IN THE NEXT CYCLE
				END IF;
			END IF;
			
			-- CHECKING CDB'S BROADCAST 
			L_0: FOR I IN 0 TO 2 LOOP 
				IF CDB_Q = RESERVATION_STATION(I)(39 DOWNTO 36) AND CDB_Q /= X"F" AND RESERVATION_STATION(I)(74) = '1' THEN -- Q RS
					RESERVATION_STATION(I)(71 DOWNTO 40) <= CDB_V; 
					RESERVATION_STATION(I)(39 DOWNTO 36) <= (OTHERS => '1'); -- Q = 1111 = VALUE IS VALID NOW
				END IF;
				IF CDB_Q = RESERVATION_STATION(I)(3 DOWNTO 0) AND CDB_Q /= X"F" AND RESERVATION_STATION(I)(74) = '1' THEN -- Q RT
					RESERVATION_STATION(I)(35 DOWNTO 4) <= CDB_V; 
					RESERVATION_STATION(I)(3 DOWNTO 0) <= (OTHERS => '1'); -- Q = 1111 = VALUE IS VALID NOW
				END IF;
			END LOOP L_0;
                        
			-- FILL RS FROM RF 
			IF RS0_WAIT_FOR_RF = '1' THEN	
				-- RS
				IF Q_RS_ROB /= "1111" THEN -- RF'S INFO IS NOT UPDATED - ROB HAS NEWER DATA
					RESERVATION_STATION(0)(71 DOWNTO 40) <= DATA_RS_ROB;
					IF DATA_RS_ROB_VALID = '1' THEN -- IS THE DATA VALID? IF YES, TAG = 1111, ELSE SAVE THE TAG GIVEN BY ROB
						RESERVATION_STATION(0)(39 DOWNTO 36) <= "1111";
					ELSE
						RESERVATION_STATION(0)(39 DOWNTO 36) <= Q_RS_ROB;
					END IF;
				ELSE -- SAVE DATA FROM RF	
					RESERVATION_STATION(0)(71 DOWNTO 40) <= DATA_RS_RF;
					RESERVATION_STATION(0)(39 DOWNTO 36) <= "1111"; --Q_RS; -- RF ALWAYS PROVIDES VALID DATA
				END IF;
				--RT
				IF Q_RT_ROB /= "1111" THEN -- RF'S INFO IS NOT UPDATED - ROB HAS NEWER DATA
					RESERVATION_STATION(0)(35 DOWNTO 4) <= DATA_RT_ROB; 
					IF DATA_RT_ROB_VALID = '1' THEN -- IS THE DATA VALID? IF YES, TAG = 1111, ELSE SAVE THE TAG GIVEN BY ROB
						RESERVATION_STATION(0)(3 DOWNTO 0) <= "1111";
					ELSE
						RESERVATION_STATION(0)(3 DOWNTO 0) <= Q_RT_ROB;
					END IF;
				ELSE -- SAVE DATA FROM RF	
					RESERVATION_STATION(0)(35 DOWNTO 4) <= DATA_RT_RF; 
					RESERVATION_STATION(0)(3 DOWNTO 0) <= "1111"; --Q_RS; -- RF ALWAYS PROVIDES VALID DATA
				END IF;
				RS0_WAIT_FOR_RF <= '0';
			ELSIF RS1_WAIT_FOR_RF = '1' THEN
				-- RS
				IF Q_RS_ROB /= "1111" THEN -- RF'S INFO IS NOT UPDATED - ROB HAS NEWER DATA
					RESERVATION_STATION(1)(71 DOWNTO 40) <= DATA_RS_ROB;
					IF DATA_RS_ROB_VALID = '1' THEN -- IS THE DATA VALID? IF YES, TAG = 1111, ELSE SAVE THE TAG GIVEN BY ROB
						RESERVATION_STATION(1)(39 DOWNTO 36) <= "1111";
					ELSE
						RESERVATION_STATION(1)(39 DOWNTO 36) <= Q_RS_ROB;
					END IF;
				ELSE -- SAVE DATA FROM RF	
					RESERVATION_STATION(1)(71 DOWNTO 40) <= DATA_RS_RF;
					RESERVATION_STATION(1)(39 DOWNTO 36) <= "1111"; --Q_RS; -- RF ALWAYS PROVIDES VALID DATA
				END IF;
				--RT
				IF Q_RT_ROB /= "1111" THEN -- RF'S INFO IS NOT UPDATED - ROB HAS NEWER DATA
					RESERVATION_STATION(1)(35 DOWNTO 4) <= DATA_RT_ROB; 
					IF DATA_RT_ROB_VALID = '1' THEN -- IS THE DATA VALID? IF YES, TAG = 1111, ELSE SAVE THE TAG GIVEN BY ROB
						RESERVATION_STATION(1)(3 DOWNTO 0) <= "1111";
					ELSE
						RESERVATION_STATION(1)(3 DOWNTO 0) <= Q_RT_ROB;
					END IF;
				ELSE -- SAVE DATA FROM RF	
					RESERVATION_STATION(1)(35 DOWNTO 4) <= DATA_RT_RF; 
					RESERVATION_STATION(1)(3 DOWNTO 0) <= "1111"; --Q_RS; -- RF ALWAYS PROVIDES VALID DATA
				END IF;
				RS1_WAIT_FOR_RF <= '0';
			ELSIF RS2_WAIT_FOR_RF = '1' THEN
				-- RS
				IF Q_RS_ROB /= "1111" THEN -- RF'S INFO IS NOT UPDATED - ROB HAS NEWER DATA
					RESERVATION_STATION(2)(71 DOWNTO 40) <= DATA_RS_ROB;
					IF DATA_RS_ROB_VALID = '1' THEN -- IS THE DATA VALID? IF YES, TAG = 1111, ELSE SAVE THE TAG GIVEN BY ROB
						RESERVATION_STATION(2)(39 DOWNTO 36) <= "1111";
					ELSE
						RESERVATION_STATION(2)(39 DOWNTO 36) <= Q_RS_ROB;
					END IF;
				ELSE -- SAVE DATA FROM RF	
					RESERVATION_STATION(2)(71 DOWNTO 40) <= DATA_RS_RF;
					RESERVATION_STATION(2)(39 DOWNTO 36) <= "1111"; --Q_RS; -- RF ALWAYS PROVIDES VALID DATA
				END IF;
				--RT
				IF Q_RT_ROB /= "1111" THEN -- RF'S INFO IS NOT UPDATED - ROB HAS NEWER DATA
					RESERVATION_STATION(2)(35 DOWNTO 4) <= DATA_RT_ROB; 
					IF DATA_RT_ROB_VALID = '1' THEN -- IS THE DATA VALID? IF YES, TAG = 1111, ELSE SAVE THE TAG GIVEN BY ROB
						RESERVATION_STATION(2)(3 DOWNTO 0) <= "1111";
					ELSE
						RESERVATION_STATION(2)(3 DOWNTO 0) <= Q_RT_ROB;
					END IF;
				ELSE -- SAVE DATA FROM RF	
					RESERVATION_STATION(2)(35 DOWNTO 4) <= DATA_RT_RF; 
					RESERVATION_STATION(2)(3 DOWNTO 0) <= "1111"; --Q_RS; -- RF ALWAYS PROVIDES VALID DATA
				END IF;
				RS2_WAIT_FOR_RF <= '0';
			END IF;
			
			-- SEND READY VALUES TO BE COMPUTED
			IF RESERVATION_STATION(0)(74) = '1' AND RESERVATION_STATION(0)(39 DOWNTO 36) = X"F" AND RESERVATION_STATION(0)(3 DOWNTO 0) = X"F" AND COUNTER < 3 THEN 
			-- IF THE RS IS BUSY AND ITS VALUES ARE READY (Q1 = Q2 = F) AND FU'S PIPELINE IS NOT FULL
				FU_Q <= RESERVATION_STATION(0)(78 DOWNTO 75); -- ROB TAG
				FU_V1 <= RESERVATION_STATION(0)(71 DOWNTO 40);
				FU_V2 <= RESERVATION_STATION(0)(35 DOWNTO 4);
				FU_OP <= RESERVATION_STATION(0)(73 DOWNTO 72);
				COUNTER <= COUNTER + 1;				
				-- RESETTING THE RS
				RESERVATION_STATION(0) <= (OTHERS => '0'); 
			ELSIF RESERVATION_STATION(1)(74) = '1' AND RESERVATION_STATION(1)(39 DOWNTO 36) = X"F" AND RESERVATION_STATION(1)(3 DOWNTO 0) = X"F" AND COUNTER < 3 THEN 
				FU_Q <= RESERVATION_STATION(1)(78 DOWNTO 75); -- ROB TAG
				FU_V1 <= RESERVATION_STATION(1)(71 DOWNTO 40);
				FU_V2 <= RESERVATION_STATION(1)(35 DOWNTO 4);
				FU_OP <= RESERVATION_STATION(1)(73 DOWNTO 72);
				COUNTER <= COUNTER + 1;
				RESERVATION_STATION(1) <= (OTHERS => '0'); 
			ELSIF RESERVATION_STATION(2)(74) = '1' AND RESERVATION_STATION(2)(39 DOWNTO 36) = X"F" AND RESERVATION_STATION(2)(3 DOWNTO 0) = X"F" AND COUNTER < 3 THEN 
				FU_Q <= RESERVATION_STATION(2)(78 DOWNTO 75); -- ROB TAG
				FU_V1 <= RESERVATION_STATION(2)(71 DOWNTO 40);
				FU_V2 <= RESERVATION_STATION(2)(35 DOWNTO 4);
				FU_OP <= RESERVATION_STATION(2)(73 DOWNTO 72);
				COUNTER <= COUNTER + 1;
				RESERVATION_STATION(2) <= (OTHERS => '0'); 
			ELSE
				FU_Q <= "1111";  -- THERE IS NO SUCH RS, WE ARE SENDING OUT NOTHING
			END IF;
			
			-- CDB JUST GOT A VALUE FROM OUR FU, UPDATING COUNTER
			IF CDB_Q_ACCESS_GRANTED = "01" AND COUNTER /= 0 THEN
				COUNTER <= COUNTER - 1;
			END IF;			
		END IF;		
	END PROCESS;
	
	ACK_SIG <= '1' WHEN (INSTRUCTION(18 DOWNTO 17) = "01" AND RST = '0' AND EXCEPTION_ROB = "1111" AND (RESERVATION_STATION(0)(74) = '0' OR RESERVATION_STATION(1)(74) = '0' OR RESERVATION_STATION(2)(74) = '0')) ELSE '0';
	ACK <= ACK_SIG;
	
END BEHAVIORAL;
