-- Computer Architecture - Technical University of Crete
-- Speculative Tomasulo’s Algorithm
-- N. Kyparissas, A. Kampylafkas

-- A DUMMY PIPELINED LOGICAL FUNCTIONAL UNIT 

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY LOGICAL_FU IS
PORT( 
	CLK 		: IN STD_LOGIC;
	RST 		: IN STD_LOGIC;
	CDB_REQ 	: OUT STD_LOGIC;
	CDB_GRANTED : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
	R1          : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	R2          : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	FOP         : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
	LOGICAL_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	Q_OUT		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	Q_IN 		: IN STD_LOGIC_VECTOR(3 DOWNTO 0));    
END LOGICAL_FU;

ARCHITECTURE BEHAVIORAL OF LOGICAL_FU IS
	TYPE Q_PIPELINE_TYPE IS ARRAY(1 DOWNTO 0) OF STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL Q_PIPELINE : Q_PIPELINE_TYPE := (OTHERS => (OTHERS => '1'));  -- "1111" THERE IS NO SUCH FU
	SIGNAL LOGICAL_RESULT_SIG 		: STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	TYPE V_PIPELINE_TYPE IS ARRAY(1 DOWNTO 0) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL V_PIPELINE : V_PIPELINE_TYPE := (OTHERS => (OTHERS => '0'));    
	SIGNAL Q_IN_SIG : STD_LOGIC_VECTOR(3 DOWNTO 0);
    
BEGIN

	LOGICAL_RESULT_SIG <= 	R1 OR R2 WHEN FOP = "00" ELSE
				R1 AND R2 WHEN FOP = "01" ELSE
				NOT R1 WHEN FOP = "10" ELSE
				(OTHERS => '0');
								
	Q_IN_SIG <= Q_IN;
	CDB_REQ <= '1' WHEN (Q_PIPELINE(1) /= "1111" AND CDB_GRANTED /= "00") OR Q_PIPELINE(0) /= "1111" ELSE '0';
	Q_OUT <= Q_PIPELINE(1);
	LOGICAL_OUT <= V_PIPELINE(1);
	
	PROCESS
	BEGIN	
		WAIT UNTIL RISING_EDGE(CLK);
		IF RST = '1' THEN
			Q_PIPELINE <= (OTHERS => (OTHERS => '1'));
		ELSE
			IF CDB_GRANTED = "00" OR Q_PIPELINE(1) = "1111" THEN
				Q_PIPELINE(1) <= Q_PIPELINE(0);
				Q_PIPELINE(0) <= Q_IN_SIG;
				V_PIPELINE(1) <= V_PIPELINE(0);
				V_PIPELINE(0) <= LOGICAL_RESULT_SIG;
			ELSIF Q_PIPELINE(0) = "1111" THEN
				Q_PIPELINE(0) <= Q_IN_SIG;
				V_PIPELINE(0) <= LOGICAL_RESULT_SIG;
 			END IF;
		END IF;
	END PROCESS;

END BEHAVIORAL;
