-- Computer Architecture - Technical University of Crete
-- Speculative Tomasulo’s Algorithm
-- N. Kyparissas, A. Kampylafkas

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;

ENTITY INSTRUCTION_FETCH IS
PORT (
	CLK : IN STD_LOGIC;
	RESET : IN STD_LOGIC;
	A_ACK : IN STD_LOGIC;
	L_ACK : IN STD_LOGIC;
	ADDR : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
	INSTRUCTION : OUT STD_LOGIC_VECTOR(18 DOWNTO 0));
END INSTRUCTION_FETCH;

ARCHITECTURE SYN OF INSTRUCTION_FETCH IS

TYPE ROM_TYPE IS ARRAY (1023 DOWNTO 0) OF STD_LOGIC_VECTOR (18 DOWNTO 0);

IMPURE FUNCTION INITROMFROMFILE (ROMFILENAME : IN STRING) RETURN ROM_TYPE IS
FILE ROMFILE : TEXT IS IN ROMFILENAME;
VARIABLE ROMFILELINE : LINE;
VARIABLE ROM : ROM_TYPE;
BEGIN
	FOR I IN 0 TO 1023 LOOP
		READLINE(ROMFILE, ROMFILELINE);
		READ (ROMFILELINE, ROM(I));
	END LOOP;
RETURN ROM;
END FUNCTION;

SIGNAL ROM : ROM_TYPE := INITROMFROMFILE("ROM.DATA");
SIGNAL ADDR_SIG : STD_LOGIC_VECTOR(9 DOWNTO 0);

BEGIN
	PROCESS
	BEGIN
	
		WAIT UNTIL RISING_EDGE(CLK);

		IF (RESET = '1') THEN
		ADDR_SIG <= (OTHERS => '0');
		ELSIF (A_ACK = '1' OR L_ACK='1') THEN 
		-- ACKS = INSTR REQUESTS COMING FROM RESERVATION STATIONS
		ADDR_SIG <= ADDR_SIG + 1;
		END IF;
			
	END PROCESS;

	INSTRUCTION <= ROM(CONV_INTEGER(ADDR_SIG));
	ADDR <= ADDR_SIG;

END SYN;


