-- Computer Architecture - Technical University of Crete
-- Speculative Tomasulo’s Algorithm
-- N. Kyparissas, A. Kampylafkas

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TOP_LEVEL IS
PORT(
	CLK : IN STD_LOGIC;
	RST : IN STD_LOGIC;
	EXCEPTION_FLAG : IN STD_LOGIC;
	EXCEPTION_ROB_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0); 
	EXCEPTION_PC : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) 
	);
END TOP_LEVEL;

ARCHITECTURE BEHAVIORAL OF TOP_LEVEL IS

	COMPONENT LOGICAL_RS_FU
	PORT(
		CLK : IN STD_LOGIC;
        RST : IN STD_LOGIC;
        -- ISSUE SIGNALS
        INSTRUCTION : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
        ACK : OUT STD_LOGIC; -- LETTING ISSUE STG KNOW THAT THIS RS IS ACCEPTING ITS CURRENT INSTR
		-- ROB SIGNALS
		Q_RS_ROB : IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- IN CASE THE DATA YOU'VE BEEN ASKING IN REGISTER FILE IS NOT VALID
		Q_RT_ROB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		DATA_RS_ROB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_RT_ROB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_RS_ROB_VALID : IN STD_LOGIC;
		DATA_RT_ROB_VALID : IN STD_LOGIC;
		Q_FOR_NEW_INSTR : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        EXCEPTION_ROB : IN STD_LOGIC_VECTOR(3 DOWNTO 0); 
		-- RF SIGNALS
		DATA_RS_RF : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_RT_RF : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		-- CDB SIGNALS
		CDB_Q : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CDB_V : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		CDB_Q_ACCESS_GRANTED : IN STD_LOGIC_VECTOR (1 DOWNTO 0); -- EVERY TIME WE SEND A VALUE TO BE COMPUTED, WE COUNT UP UNTIL THE PIPELINE IS FULL.
											-- EVERY TIME CDB TAKES A VALUE, WE COUNT DOWN AND THAT MEANS WE CAN SEND ANOTHER VALUE. 
		CDB_REQ 		: OUT STD_LOGIC;
		LOGICAL_OUT  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		Q_OUT			: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
	END COMPONENT;

	COMPONENT ARITHMETIC_RS_FU
    PORT(
        CLK : IN STD_LOGIC;
        RST : IN STD_LOGIC;
        -- ISSUE SIGNALS
        INSTRUCTION : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
        ACK : OUT STD_LOGIC; -- LETTING ISSUE STG KNOW THAT THIS RS IS ACCEPTING ITS CURRENT INSTR
		-- ROB SIGNALS
		Q_RS_ROB : IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- IN CASE THE DATA YOU'VE BEEN ASKING IN REGISTER FILE IS NOT VALID
		Q_RT_ROB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		DATA_RS_ROB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_RT_ROB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_RS_ROB_VALID : IN STD_LOGIC;
		DATA_RT_ROB_VALID : IN STD_LOGIC;
		Q_FOR_NEW_INSTR : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        EXCEPTION_ROB : IN STD_LOGIC_VECTOR(3 DOWNTO 0); 
		-- RF SIGNALS
		DATA_RS_RF : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_RT_RF : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        -- CDB SIGNALS
        CDB_Q : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        CDB_V : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        CDB_Q_ACCESS_GRANTED : IN STD_LOGIC_VECTOR (1 DOWNTO 0); -- EVERY TIME WE SEND A VALUE TO BE COMPUTED, WE COUNT UP UNTIL THE PIPELINE IS FULL.
                                            -- EVERY TIME CDB TAKES A VALUE, WE COUNT DOWN AND THAT MEANS WE CAN SEND ANOTHER VALUE. 
        CDB_REQ 		: OUT STD_LOGIC;
        ARITHMETIC_OUT  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        Q_OUT			: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
	END COMPONENT;

	COMPONENT INSTRUCTION_FETCH
    PORT( 
        A_ACK       : IN STD_LOGIC;
        L_ACK       : IN STD_LOGIC;
        RESET		: IN STD_LOGIC;
        ADDR 		: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
        CLK  		: IN STD_LOGIC;
        INSTRUCTION : OUT STD_LOGIC_VECTOR(18 DOWNTO 0));
	END COMPONENT;

	COMPONENT CDB
    PORT ( 
           ARITHMETIC_REQ : IN STD_LOGIC;
           LOGICAL_REQ : IN STD_LOGIC;
           ARITHMETIC_DATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
           LOGICAL_DATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
           ARD_Q : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
           LRD_Q : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
           CLK : IN STD_LOGIC;
           RESET : IN STD_LOGIC;
           GRANTED : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
           CDB_VALUE : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
           CDB_Q : OUT STD_LOGIC_VECTOR (3 DOWNTO 0));
	END COMPONENT;

	COMPONENT REGISTER_FILE
    PORT( 
		CLK : IN STD_LOGIC;
		RST : IN STD_LOGIC;
		-- ROB
		ROB_RD : IN STD_LOGIC_VECTOR(4 DOWNTO 0); 
		ROB_V : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		ROB_WE : IN STD_LOGIC;
		-- RF PORTS
		RS : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		RT : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		DATA_RS : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_RT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
	END COMPONENT;

	COMPONENT ROB 
	PORT (
		CLK : IN STD_LOGIC;
		RST : IN STD_LOGIC;
		-- ISSUE
		PC : IN STD_LOGIC_VECTOR(9 DOWNTO 0); -- HERE: OUR PC COUNTER
		ISSUE_WE : IN STD_LOGIC;
		INSTRUCTION : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
		Q_FOR_NEW_INSTR : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); -- = TAIL 
		-- NEW INSTRUCTION
		Q_RS_ROB : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); -- IN CASE THE DATA YOU'VE BEEN ASKING IN REGISTER FILE IS NOT VALID
		Q_RT_ROB : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		DATA_RS_ROB : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_RT_ROB : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_RS_ROB_VALID : OUT STD_LOGIC;
		DATA_RT_ROB_VALID : OUT STD_LOGIC;
		-- CDB
		CDB_V : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		CDB_Q : IN STD_LOGIC_VECTOR(3 DOWNTO 0); 
		-- RF (COMMIT)
		ROB_VALUE : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		ROB_RD : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		RF_WE : OUT STD_LOGIC;
		-- EXCEPTION
		EXCEPTION_PC : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		EXCEPTION_ROB_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); -- NOTIFYING RS WHICH ROBS TO FLUSH 
		EXCEPTION_FLAG : IN STD_LOGIC; 
		EXCEPTION_ROB_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0));
	END COMPONENT;

	SIGNAL A_ACK, L_ACK, ISSUE_WE, CDB_REQ_L, CDB_REQ_A, RF_WE, DATA_RS_ROB_VALID, DATA_RT_ROB_VALID: STD_LOGIC := '0';
	SIGNAL INSTRUCTION : STD_LOGIC_VECTOR(18 DOWNTO 0) := (OTHERS => '1');
	SIGNAL CDB_Q, Q_FOR_NEW_INSTR, Q_RS_ROB, Q_RT_ROB, Q_L, Q_A, EXCEPTION_ROB_OUT : STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '1'); 
	SIGNAL CDB_V, DATA_RS_RF, DATA_RT_RF, DATA_RS_ROB, DATA_RT_ROB, ROB_V, ARITHMETIC_DATA, LOGICAL_DATA : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0'); 
	SIGNAL CDB_Q_ACCESS_GRANTED : STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '1'); 
	SIGNAL PC : STD_LOGIC_VECTOR(9 DOWNTO 0) := (OTHERS => '0');
	SIGNAL ROB_RD : STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
	
BEGIN

	ISSUE_CP: INSTRUCTION_FETCH
	PORT MAP(   
		A_ACK => A_ACK,
		L_ACK => L_ACK,
		RESET  => RST,
		CLK   => CLK,
		ADDR => PC,
		INSTRUCTION => INSTRUCTION);

	ISSUE_WE <= A_ACK OR L_ACK;

	RF: REGISTER_FILE
	PORT MAP( 
		CLK => CLK,
		RST => RST,
		ROB_RD => ROB_RD, 
		ROB_V => ROB_V,
		ROB_WE => RF_WE,
		RS => INSTRUCTION(9 DOWNTO 5),
		RT => INSTRUCTION(4 DOWNTO 0),
		DATA_RS => DATA_RS_RF, 
		DATA_RT => DATA_RT_RF);

	LRS: LOGICAL_RS_FU
	PORT MAP(
		CLK => CLK,
		RST => RST,
		INSTRUCTION => INSTRUCTION,
		ACK => L_ACK,
		-- ROB SIGNALS
		Q_RS_ROB => Q_RS_ROB,
		Q_RT_ROB => Q_RT_ROB,
		DATA_RS_ROB => DATA_RS_ROB,
		DATA_RT_ROB => DATA_RT_ROB,
		DATA_RS_ROB_VALID => DATA_RS_ROB_VALID,
		DATA_RT_ROB_VALID => DATA_RT_ROB_VALID,
		Q_FOR_NEW_INSTR => Q_FOR_NEW_INSTR,
        EXCEPTION_ROB => EXCEPTION_ROB_OUT,
		-- RF SIGNALS
		DATA_RS_RF => DATA_RS_RF,
		DATA_RT_RF => DATA_RT_RF,
		-- CDB SIGNALS
		CDB_Q => CDB_Q,
		CDB_V => CDB_V,
		CDB_Q_ACCESS_GRANTED => CDB_Q_ACCESS_GRANTED,
		CDB_REQ => CDB_REQ_L,
		LOGICAL_OUT => LOGICAL_DATA,
		Q_OUT => Q_L);

	ARS: ARITHMETIC_RS_FU
	PORT MAP(
		CLK => CLK,
		RST => RST,
		INSTRUCTION => INSTRUCTION,
		ACK => A_ACK,
		-- ROB SIGNALS
		Q_RS_ROB => Q_RS_ROB,
		Q_RT_ROB => Q_RT_ROB,
		DATA_RS_ROB => DATA_RS_ROB,
		DATA_RT_ROB => DATA_RT_ROB,
		DATA_RS_ROB_VALID => DATA_RS_ROB_VALID,
		DATA_RT_ROB_VALID => DATA_RT_ROB_VALID,
		Q_FOR_NEW_INSTR => Q_FOR_NEW_INSTR,
        EXCEPTION_ROB => EXCEPTION_ROB_OUT,
		-- RF SIGNALS
		DATA_RS_RF => DATA_RS_RF,
		DATA_RT_RF => DATA_RT_RF,
		-- CDB SIGNALS
		CDB_Q => CDB_Q,
		CDB_V => CDB_V,
		CDB_Q_ACCESS_GRANTED => CDB_Q_ACCESS_GRANTED,
		CDB_REQ => CDB_REQ_A,
		ARITHMETIC_OUT => ARITHMETIC_DATA,
		Q_OUT => Q_A);

	CDBS: CDB
	PORT MAP( 
		ARITHMETIC_REQ => CDB_REQ_A,
		LOGICAL_REQ => CDB_REQ_L,
		ARITHMETIC_DATA => ARITHMETIC_DATA,
		LOGICAL_DATA => LOGICAL_DATA,
		ARD_Q => Q_A,
		LRD_Q => Q_L,
		CLK => CLK,
		RESET => RST,
		GRANTED => CDB_Q_ACCESS_GRANTED,
		CDB_VALUE => CDB_V,
		CDB_Q => CDB_Q);
		   
	ROBBING_IN_ORDER: ROB
	PORT MAP(
		CLK => CLK,
		RST => RST,
		-- ISSUE
		PC => PC,
		ISSUE_WE => ISSUE_WE,
		INSTRUCTION => INSTRUCTION,
		-- ROB SIGNALS
		Q_RS_ROB => Q_RS_ROB,
		Q_RT_ROB => Q_RT_ROB,
		DATA_RS_ROB => DATA_RS_ROB,
		DATA_RT_ROB => DATA_RT_ROB,
		DATA_RS_ROB_VALID => DATA_RS_ROB_VALID,
		DATA_RT_ROB_VALID => DATA_RT_ROB_VALID,
		Q_FOR_NEW_INSTR => Q_FOR_NEW_INSTR,
		-- CDB
		CDB_V => CDB_V,
		CDB_Q => CDB_Q,
		-- RF (COMMIT)
		ROB_VALUE => ROB_V,
		ROB_RD => ROB_RD,
		RF_WE => RF_WE,
		-- EXCEPTION
		EXCEPTION_PC => EXCEPTION_PC,
		EXCEPTION_ROB_OUT => EXCEPTION_ROB_OUT,
		EXCEPTION_FLAG => EXCEPTION_FLAG,
		EXCEPTION_ROB_IN => EXCEPTION_ROB_IN);

END BEHAVIORAL;
