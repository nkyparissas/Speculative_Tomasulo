-- Computer Architecture - Technical University of Crete
-- Speculative Tomasulo’s Algorithm
-- N. Kyparissas, A. Kampylafkas

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY CDB IS 
PORT ( 
	ARITHMETIC_REQ : IN STD_LOGIC;
	LOGICAL_REQ : IN STD_LOGIC;
	ARITHMETIC_DATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	LOGICAL_DATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	ARD_Q : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	LRD_Q : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	CLK : IN STD_LOGIC;
	RESET : IN STD_LOGIC;
	GRANTED : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
	CDB_VALUE : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
	CDB_Q : OUT STD_LOGIC_VECTOR (3 DOWNTO 0));
END CDB;

ARCHITECTURE BEHAVIORAL OF CDB IS
    SIGNAL PREV : STD_LOGIC_VECTOR (1 DOWNTO 0) := "01";
    SIGNAL CDB_GRANTED, OUTPUT_SEL : STD_LOGIC_VECTOR (1 DOWNTO 0) := "11";
 
BEGIN

    PROCESS
    BEGIN
        WAIT UNTIL(CLK'EVENT AND CLK = '1');
        
        IF(RESET='1')THEN
            CDB_GRANTED <= "11"; -- "11" MEANS NO ONE GETS ACCESS TO CDB
            PREV <= "01";		 -- INITIALIZING PRIORITY TO LOGICAL / SUPPOSING ARITHMETIC WAS THE PREVIOUS ONE TO ACCESS CDB
		-- BOTH REQUEST ACCESS TO CDB, SO WE CHECK WHO HAD ACCESS THE PREVIOUS TIME	
        ELSIF(ARITHMETIC_REQ = '1' AND LOGICAL_REQ = '1')THEN
            IF(PREV="01")THEN -- GRANTING ACCESS TO LOGICAL
                CDB_GRANTED <= "00";
                PREV <= "00";		
            ELSE
                CDB_GRANTED <= "01";
                PREV <= "01";	
            END IF;
        ELSIF(ARITHMETIC_REQ = '1')THEN
            CDB_GRANTED <= "01";
            PREV <= "01";		
        ELSIF(LOGICAL_REQ = '1')THEN
            CDB_GRANTED <= "00";
            PREV <= "00";		
        ELSE       
            CDB_GRANTED <= "11";
        END IF;        
        
    END PROCESS;
	
	OUTPUT_SEL <= CDB_GRANTED;
	
	GRANTED <= CDB_GRANTED;
	
	CDB_VALUE <= 	ARITHMETIC_DATA WHEN OUTPUT_SEL = "01" ELSE
					LOGICAL_DATA WHEN OUTPUT_SEL = "00" ELSE
					(OTHERS => '0');
				
	CDB_Q <=    ARD_Q WHEN OUTPUT_SEL = "01" ELSE
				LRD_Q WHEN OUTPUT_SEL = "00" ELSE
				(OTHERS => '1');
				
END BEHAVIORAL;
