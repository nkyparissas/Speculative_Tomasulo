-- Computer Architecture - Technical University of Crete
-- Speculative Tomasulo’s Algorithm
-- N. Kyparissas, A. Kampylafkas

-- TESTBENCH AUTOMATICALLY GENERATED ONLINE
-- AT HTTP://VHDL.LAPINOO.NET
-- GENERATION DATE : 13.12.2017 15:21:11 GMT

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TB_TOP_LEVEL IS
END TB_TOP_LEVEL;

ARCHITECTURE TB OF TB_TOP_LEVEL IS

	COMPONENT TOP_LEVEL
	PORT (
		CLK              : IN STD_LOGIC;
		RST              : IN STD_LOGIC;
		EXCEPTION_FLAG   : IN STD_LOGIC;
		EXCEPTION_ROB_IN : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		EXCEPTION_PC     : OUT STD_LOGIC_VECTOR (9 DOWNTO 0));
	END COMPONENT;

	SIGNAL CLK              : STD_LOGIC;
	SIGNAL RST              : STD_LOGIC;
	SIGNAL EXCEPTION_FLAG   : STD_LOGIC;
	SIGNAL EXCEPTION_ROB_IN : STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL EXCEPTION_PC     : STD_LOGIC_VECTOR (9 DOWNTO 0);

	CONSTANT TBPERIOD : TIME := 10 NS; 
	SIGNAL TBCLOCK : STD_LOGIC := '1';
	SIGNAL TBSIMENDED : STD_LOGIC := '0';

BEGIN

	DUT : TOP_LEVEL
	PORT MAP (
		CLK              => CLK,
		RST              => RST,
		EXCEPTION_FLAG   => EXCEPTION_FLAG,
		EXCEPTION_ROB_IN => EXCEPTION_ROB_IN,
		EXCEPTION_PC     => EXCEPTION_PC);

    -- CLOCK GENERATION
    TBCLOCK <= NOT TBCLOCK AFTER TBPERIOD/2 WHEN TBSIMENDED /= '1' ELSE '0';

    -- EDIT: CHECK THAT CLK IS REALLY YOUR MAIN CLOCK SIGNAL
    CLK <= TBCLOCK;

    STIMULI : PROCESS
    BEGIN
        -- EDIT ADAPT INITIALIZATION AS NEEDED
        EXCEPTION_FLAG <= '0';
        EXCEPTION_ROB_IN <= (OTHERS => '0');

        -- RESET GENERATION
        -- EDIT: CHECK THAT RST IS REALLY YOUR RESET SIGNAL
        RST <= '1';
        WAIT FOR 2 * TBPERIOD;
        RST <= '0';
        WAIT FOR 1 * TBPERIOD;
        
        -- -- EXCEPTION
        -- -- ROB 0 - 4 FULL, EXCEPTION AT ROB 3 
        -- -- MUST FLUSH: ROB 3 + ROB 4, RS_LOGICAL[0] + RS_ARITH[1]
         WAIT FOR 5 * TBPERIOD;
         EXCEPTION_FLAG <= '1';
         EXCEPTION_ROB_IN <= "0011";
         WAIT FOR 1 * TBPERIOD;
         EXCEPTION_FLAG <= '0';
        -- -- END OF EXCEPTION
        
        -- EDIT ADD STIMULI HERE
        WAIT FOR 100 * TBPERIOD;

        -- STOP THE CLOCK AND HENCE TERMINATE THE SIMULATION
        TBSIMENDED <= '1';
        WAIT;
    END PROCESS;

END TB;