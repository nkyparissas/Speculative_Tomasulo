-- Computer Architecture - Technical University of Crete
-- Speculative Tomasulo’s Algorithm
-- N. Kyparissas, A. Kampylafkas

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ARITHMETIC_RS_FU IS
PORT(
	CLK : IN STD_LOGIC;
	RST : IN STD_LOGIC;
	-- ISSUE SIGNALS
	INSTRUCTION : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
	ACK : OUT STD_LOGIC; -- LETTING ISSUE STG KNOW THAT THIS RS IS ACCEPTING ITS CURRENT INSTR
	-- ROB SIGNALS
	Q_RS_ROB : IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- IN CASE THE DATA YOU'VE BEEN ASKING IN REGISTER FILE IS NOT VALID
	Q_RT_ROB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	DATA_RS_ROB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	DATA_RT_ROB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	DATA_RS_ROB_VALID : IN STD_LOGIC;
	DATA_RT_ROB_VALID : IN STD_LOGIC;
	Q_FOR_NEW_INSTR : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	EXCEPTION_ROB : IN STD_LOGIC_VECTOR(3 DOWNTO 0); 
	-- RF SIGNALS
	DATA_RS_RF : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	DATA_RT_RF : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	-- CDB SIGNALS
	CDB_Q : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	CDB_V : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	CDB_Q_ACCESS_GRANTED : IN STD_LOGIC_VECTOR (1 DOWNTO 0); -- EVERY TIME WE SEND A VALUE TO BE COMPUTED, WE COUNT UP UNTIL THE PIPELINE IS FULL.
										-- EVERY TIME CDB TAKES A VALUE, WE COUNT DOWN AND THAT MEANS WE CAN SEND ANOTHER VALUE. 
	CDB_REQ 		: OUT STD_LOGIC;
	ARITHMETIC_OUT  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	Q_OUT			: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END ARITHMETIC_RS_FU;

ARCHITECTURE BEHAVIORAL OF ARITHMETIC_RS_FU IS
    SIGNAL FU_OP : STD_LOGIC_VECTOR(1 DOWNTO 0);
    SIGNAL FU_Q : STD_LOGIC_VECTOR(3 DOWNTO 0);     
    SIGNAL FU_V1, FU_V2 : STD_LOGIC_VECTOR(31 DOWNTO 0);

    COMPONENT RESERVATION_STATIONS_ARITH 
	PORT(
		CLK : IN STD_LOGIC;
		RST : IN STD_LOGIC;
		-- ISSUE SIGNALS
		INSTRUCTION : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
		ACK : OUT STD_LOGIC; -- LETTING ISSUE STG KNOW THAT THIS RS IS ACCEPTING ITS CURRENT INSTR
		-- ROB SIGNALS
		Q_RS_ROB : IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- IN CASE THE DATA YOU'VE BEEN ASKING IN REGISTER FILE IS NOT VALID
		Q_RT_ROB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		DATA_RS_ROB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_RT_ROB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_RS_ROB_VALID : IN STD_LOGIC;
		DATA_RT_ROB_VALID : IN STD_LOGIC;
		Q_FOR_NEW_INSTR : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		EXCEPTION_ROB : IN STD_LOGIC_VECTOR(3 DOWNTO 0); 
		-- RF SIGNALS
		DATA_RS_RF : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_RT_RF : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		-- FU SIGNALS
		FU_Q : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);  
		FU_V1 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		FU_V2 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		FU_OP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		-- CDB SIGNALS
		CDB_Q : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CDB_V : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		CDB_Q_ACCESS_GRANTED : IN STD_LOGIC_VECTOR (1 DOWNTO 0)); 
    END COMPONENT;

    COMPONENT ARITHMETIC_FU 
	PORT( 
		CLK 			: IN STD_LOGIC;
		RST 			: IN STD_LOGIC;
		CDB_REQ 		: OUT STD_LOGIC;
		CDB_GRANTED		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		R1              : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		R2              : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		FOP             : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		ARITHMETIC_OUT  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		Q_OUT			: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		Q_IN            : IN STD_LOGIC_VECTOR(3 DOWNTO 0));      
    END COMPONENT;

BEGIN

	RS: RESERVATION_STATIONS_ARITH 
    PORT MAP(
		CLK => CLK,
		RST => RST,
		-- ISSUE SIGNALS
		INSTRUCTION => INSTRUCTION,
		ACK => ACK, 
		-- ROB SIGNALS
		Q_RS_ROB => Q_RS_ROB,
		Q_RT_ROB => Q_RT_ROB,
		DATA_RS_ROB => DATA_RS_ROB,
		DATA_RT_ROB => DATA_RT_ROB,
		DATA_RS_ROB_VALID => DATA_RS_ROB_VALID,
		DATA_RT_ROB_VALID => DATA_RT_ROB_VALID,
		Q_FOR_NEW_INSTR => Q_FOR_NEW_INSTR,
		EXCEPTION_ROB => EXCEPTION_ROB,
		-- RF SIGNALS
		DATA_RS_RF => DATA_RS_RF,
		DATA_RT_RF => DATA_RT_RF,
		-- INTERNAL SIGNALS
		FU_Q => FU_Q,  
		FU_V1 => FU_V1,
		FU_V2 => FU_V2,
		FU_OP => FU_OP,
		-------------------
		CDB_Q => CDB_Q,
		CDB_V => CDB_V,
		CDB_Q_ACCESS_GRANTED => CDB_Q_ACCESS_GRANTED);

	FU: ARITHMETIC_FU 
    PORT MAP( 
        CLK => CLK,
		RST => RST,
		CDB_REQ => CDB_REQ,
		CDB_GRANTED => CDB_Q_ACCESS_GRANTED,
		-- INTERNAL SIGNALS
		R1 => FU_V1,
        R2 => FU_V2,
        FOP => FU_OP,
        Q_IN => FU_Q,
        -------------------
        ARITHMETIC_OUT  => ARITHMETIC_OUT,
		Q_OUT => Q_OUT);  

END BEHAVIORAL;